/* -------------------------------------------------------------  
   COMBINATIONAL CIRCUIT | OR GATE
---------------------------------------------------------------- */

module or_gate
(
	input a,
	input b,
	output y
);
assign y = a | b;
endmodule

/* -------------------------------------------------------------  
                        2024 NIGIL M R
---------------------------------------------------------------- */